module ID(instruction, opcode, Rn, Rm, Rd, funct7, funct3, imm12, );



endmodule
