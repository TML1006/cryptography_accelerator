module forwardingLogic();
	//If instruction in mem mix columns stage shares register send the output ahead and mux with the old value
	//Any spot before that should also receive if it is in reg/dec stage
	
	
	//Same for encryption forward the appropriate value
	
	


endmodule
